library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

use work.common_pack.all;

library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

entity cmdProc is
port(
 clk:		in std_logic;
 reset:		in std_logic;
 rxnow:		in std_logic;
 rxData:    in std_logic_vector (7 downto 0);
 txData:	out std_logic_vector (7 downto 0);
 rxdone:	out std_logic;
 ovErr:		in std_logic;
 framErr:	in std_logic;
 txnow:		out std_logic;
 txdone:	in std_logic;
 start:     out std_logic;
 numWords_bcd:out BCD_ARRAY_TYPE(2 downto 0);
 dataReady: in std_logic;
 byte:      in std_logic_vector(7 downto 0);
 maxIndex:  in BCD_ARRAY_TYPE(2 downto 0);
 dataResults:in CHAR_ARRAY_TYPE(0 to RESULT_BYTE_NUM-1);
 seqDone:   in std_logic
  );
end;

ARCHITECTURE myarch OF cmdProc IS

  COMPONENT counter
	PORT (
     clk: in std_logic;
     rst: in std_logic;
     en: in std_logic;
     cntOut: out std_logic_vector(5 downto 0)
     );
     END COMPONENT;
     SIGNAL rst0, en0:STD_LOGIC; 
     SIGNAL cnt0Out:STD_LOGIC_VECTOR(5 downto 0);

  COMPONENT reg
    PORT (
	 clk: in std_logic;
	 regreset: in std_logic;
     load: in std_logic;
     D: in std_logic_vector(7 downto 0);
     Q: out std_logic_vector(7 downto 0)
     );
     END COMPONENT;
     SIGNAL regreset0, load0: std_logic;
     SIGNAL D0, Q0: std_logic_vector(7 downto 0);
	
  COMPONENT shift
	 PORT (
      shift_in : in std_logic_vector(7 downto 0); -- DATA IN
      en_shift : in std_logic; -- CHIP ENABLE
      load_shift : in std_logic;
      clk : in std_logic; -- CLOCK
      shift_out : out BCD_ARRAY_TYPE(2 downto 0) -- SHIFTER OUTPUT
      );
      END COMPONENT;
      SIGNAL shift_in: std_logic_vector(7 downto 0);              
      SIGNAL shift_out: BCD_ARRAY_TYPE(2 downto 0);
      SIGNAL en1, load1 : std_logic;
      
  COMPONENT seqdonecounter
    PORT(
     clk : in std_logic;
     rst : in std_logic;
     en : in std_logic;
     SEQcntOut : out std_logic_vector(1 downto 0)
     );
     END COMPONENT;
     SIGNAL rst_SeqDone, en_SeqDone:STD_LOGIC; 
     SIGNAL SEQcntOut:STD_LOGIC_VECTOR(1 downto 0);
      
  COMPONENT byteMux
     PORT ( 
      clk : in std_logic;
      data : in std_logic_vector(3 downto 0);
      address : in std_logic_vector(5 downto 0);
      q: out  std_logic_vector(7 downto 0)
      );
      END COMPONENT;   
      SIGNAL data: std_logic_vector(3 downto 0);
      SIGNAL address: std_logic_vector(5 downto 0);   
      SIGNAL q: std_logic_vector(7 downto 0);
      
  COMPONENT formatmux is
    PORT ( 
        clk : in std_logic;
        countIn : in std_logic_vector(5 downto 0);
        formatout: out std_logic_vector(7 downto 0)
        );
        END COMPONENT; 
        SIGNAL countIn: std_logic_vector(5 downto 0);   
        SIGNAL formatout: std_logic_vector(7 downto 0);
     
     
  FOR cnt0: counter USE ENTITY work.myCounter(Behavioral); 
  FOR reg0: reg USE ENTITY work.myRegister(Behavioral);
  FOR shift0: shift USE ENTITY work.shift(shift_arch);  
  FOR Seqcnt: seqdonecounter USE ENTITY work.seqdonecounter(Behavioral);
  FOR mux1: bytemux USE ENTITY work.bytemux(mux);
  FOR mux2: formatmux USE ENTITY work.formatmux(Behavioral);
 
  TYPE state_type IS (STATE1, INIT, COUNT_CHECK, A_CHECK, NUM_CHECK, ERROR, CORRECT_WORD, 
  SHIFTER, WAIT_SHIFT, FORMAT1, FORMAT2, FORMAT3, WAIT_FORMAT, FORMAT_CHECK, SEQ_CHECK, FINAL_FORMAT, START1, DATA_WAIT,WAIT_BYTE,
  LOAD_BYTE, LAST_BYTE, BYTE1, TRANSMIT1, WAIT_TX, LOAD_BYTE2, BYTE2, TRANSMIT2, WAIT_TX2 ); 
  SIGNAL curState, nextState: state_type;


BEGIN 
 cnt0: counter PORT MAP(clk, rst0, en0, cnt0Out);
 reg0: reg PORT MAP(clk, regreset0, load0, D0, Q0); 
 shift0: shift PORT MAP(shift_in,en1,load1,clk,shift_out);
 Seqcnt: SeqDoneCounter PORT MAP(clk,rst_SeqDone,en_SeqDone,SEQcntOut);
 mux1: ByteMUX PORT MAP(clk,data,address,q);
 mux2: formatmux PORT MAP(clk,countIn,formatout);
 
 combi_nextState: PROCESS(curState, rxNow, rxData, cnt0Out,txdone,dataready,SEQcntOut)
  BEGIN    
    CASE curState IS
	
	WHEN STATE1 =>
	nextState <= INIT;
	
	WHEN INIT =>
	 if rxNow = '1' then 
		nextState <= COUNT_CHECK;
	 else 
		nextState <= curState;
	 end if; 
	 
	WHEN COUNT_CHECK =>
	 if cnt0Out = "000000" then
	    nextState <= A_CHECK;
	 else
		nextState <= NUM_CHECK;
	 end if;
	 
	WHEN A_CHECK =>
	 if rxData = "01000001" then --if dataIn = A
	    nextState <= CORRECT_WORD;
	 elsif rxData = "01100001" then --if dataIn = a
	    nextState <= CORRECT_WORD;
	 else
		nextState<= ERROR;
	 end if;
	 
	WHEN NUM_CHECK =>
	 if (rxData >= "00110000") and (rxData <= "00111001") then  --0
		nextState <= CORRECT_WORD;
	else 
		nextState <= ERROR;
	end if; 
	
	WHEN ERROR => 
     nextState <= curState;
	  
	WHEN CORRECT_WORD =>
	  if (cnt0Out <= "000011") and (cnt0Out > "000000" ) then
	  nextState <= SHIFTER;                                 
	  elsif 
      cnt0Out = "000000" then 
      nextState <= INIT;
	  else
	  nextState <= curState;
	  end if; 
 
   WHEN SHIFTER =>
	 if cnt0Out >= "000100"  then 
	 NextState <= WAIT_SHIFT;        
	 else  
	   nextState <= INIT;
	 end if;
	
	WHEN WAIT_SHIFT =>
	 if txdone ='1' then
	  nextState <= FORMAT1;
    else
	  nextState <= curState;
	  end if; 
	  
	WHEN FORMAT1 =>
	  nextState <= FORMAT2;
	
	WHEN FORMAT2 =>
	  nextState <= FORMAT3;
	   
	WHEN FORMAT3 =>         
	   nextState <= WAIT_FORMAT;
    
    WHEN WAIT_FORMAT =>
       if txdone = '1' then 
       nextState <= FORMAT_CHECK;
       else    
	   nextState <= curState; 
	   end if;
	
	WHEN FORMAT_CHECK =>
	  if cnt0Out > "001001" then
	   nextState <= SEQ_CHECK;
	   else
	   nextState <= FORMAT1;
	   end if; 
	
	WHEN SEQ_CHECK =>    
	  if SEQcntOut = "01" then
	    nextState <= FINAL_FORMAT;
	  elsif SEQcntOut = "10" then
	    nextState <= STATE1;
	  else 
	    nextState <= START1; 
	  end if;                 
	
	WHEN FINAL_FORMAT =>
	   nextState <= FORMAT1;
	
	WHEN START1 =>
	  nextState <= DATA_WAIT; 
	
	WHEN DATA_WAIT =>
	  if dataready = '1' then
	  nextState <= WAIT_BYTE;
	  else 
	  nextState <= CurState;
   	  end if;
   	
   	WHEN WAIT_BYTE =>   
   	  nextState <= LOAD_BYTE;
   	  
   	WHEN LOAD_BYTE =>
   	  if seqDone = '1' then
	  nextState <= LAST_BYTE; 
	  else
   	  nextState <= BYTE1;
   	  end if;
   	
   	WHEN LAST_BYTE =>
   	  nextState <= TRANSMIT1;
   	
   	WHEN BYTE1 =>
	  nextState <= TRANSMIT1;
	  
	WHEN TRANSMIT1 =>
	  nextState <= WAIT_TX; 
          	
	WHEN WAIT_TX =>
	  if txDone = '1' then      
 	    nextState <= LOAD_BYTE2;
	  else
	    nextState <= curState;
	  end if; 
	
	WHEN LOAD_BYTE2 =>
	  nextState <= BYTE2;
	
	WHEN BYTE2 =>
	  nextState <= TRANSMIT2; 
	  
	WHEN TRANSMIT2 =>      
	   nextState <= WAIT_TX2; 
	
	WHEN WAIT_TX2 =>
	  if txDone = '1' then      
 	    nextState <= FORMAT1;
	  else
	    nextState <= curState;
	  end if; 
	 
	 WHEN others =>
	   nextState <= INIT;
	
    end CASE;
  end PROCESS; 

  combi_out: PROCESS(curState)
  BEGIN
  
  --inital conditions 
  D0 <= "00000000"; 
  en0 <= '0';
  rst0 <= '0';
  regreset0 <= '0';
  load0 <= '0';
  load1 <= '0';
  rxdone <= '0';
  txData <= Q0;
  txnow <= '0';
  en1 <= '0';
  shift_in <= rxdata;
  start <= '0';
  numWords_bcd <= shift_out;
  address <= cnt0Out;
  en_SeqDone <= '0';
  rst_SeqDone <= '0';
  countIn <= cnt0Out;
  --if curState = INIT then 
  --INITIAL CONDITIONS 
  --end if;
  if curState = STATE1 then
  rst0 <= '1';
  rst_SeqDone <= '1';
  end if;
  
  if curState = COUNT_CHECK then
  D0 <= rxData;
  load0 <= '1';
  end if;
  
  if curState = A_CHECK then 
  txnow <= '1';
  end if; 
  
  if curState = NUM_CHECK then 
  txnow <= '1'; 
  end if; 
  
  if curState = ERROR then 
  rst0 <= '1';
  rxdone <= '1';
    end if; 
  
  if curState = CORRECT_WORD then 
  en0 <= '1';
  rxdone <= '1';-- need to find number of clock cycles for when there are 3 numbers. 
    end if; 
  
  if curState = SHIFTER then
  en1 <= '1';
  end if;

  if curState = WAIT_SHIFT then 
  load1 <= '1'; 
  --NNN
  end if; 
  
  if curState = FORMAT1 then
  en0 <= '1';
  D0 <= formatout;
  load0 <= '1';
  END IF;
                                   
  if curState = FORMAT2 then
    END IF;
  
  if curState = FORMAT3 then               
  txnow <= '1';              
  END IF;    
                  
  if curState = FINAL_FORMAT then
  rst0 <= '1';
  en_SeqDone <= '1';
  end if;
  
  if curState = START1 then  
  start <= '1';            
  end if; 
  
  if curState = DATA_WAIT then
  end if;
  
  if curState = WAIT_BYTE then
  data <= byte(7 downto 4);
  
  end if;
  
  if curState = LAST_BYTE then
  en_SeqDone <= '1';
  end if;
  
  if curState = LOAD_BYTE then
  D0 <= q;
  load0 <= '1';
  end if;
  
  if curState = BYTE1 then 
   end if; 
  
  if curState = TRANSMIT1 then
  txnow <= '1';
  en0 <= '1';
  end if;                 
  
  if curState = WAIT_TX then
  data <= byte(3 downto 0);
  end if;
  
  if curState = LOAD_BYTE2 then
  D0 <= q;
  load0 <= '1';
  end if;
  
  if curState = BYTE2 then
  end if;      
  
  if curState = TRANSMIT2 then
  txnow <= '1';
  end if;                                
                              
  END PROCESS; 

  seq_state: PROCESS (clk, reset)
  BEGIN
    if reset = '1' then
      curState <= STATE1;
    elsif clk'EVENT AND clk='1' then
      curState <= nextState;
    end if;
  end PROCESS;
end;